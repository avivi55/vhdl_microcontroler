library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_signed.all;

entity microcontroller is
    port (
        clock : in std_logic
    );
end entity;